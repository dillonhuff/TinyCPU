module write_detector(input [31:0] instruction,

                      output       writes_reg,
                      output [4:0] register);

   
endmodule
