module RAW_dependence_detector(input [31:0] );
   
endmodule
