module cpu();

   
endmodule
