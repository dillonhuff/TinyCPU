module cpu_pipelined_basic();
endmodule
