module stall_detector(output [0:0] stall);

   assign stall = 1'b0;

endmodule
