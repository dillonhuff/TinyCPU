module stage_decode();
endmodule
