module read_detector(input [31:0] instr,
                     
                     output reads_0,
                     output reads_1,

                     output [4:0] read_reg_0,
                     output [4:0] read_reg_1);
endmodule
