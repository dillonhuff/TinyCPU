module decoder();


endmodule
